
library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;
use work.video_stream_pkg.all;

entity VIDEO_PROCESSING is
generic(W : integer := 16);
    port(
        clk       		: in  std_logic;
        sresetn   		: in  std_logic;
        videoStreamIn   : in  VideoStream_t;
		AUDIO_IN		: in std_logic_vector(W-1 downto 0);
        videoStreamOut  : out VideoStream_t
    );

end entity;

architecture RTL of VIDEO_PROCESSING is

-- video parameters ----------------------------------
	-- screen size in pixels incl. blank region
	constant X_FULL : natural := 1040; 
	constant Y_FULL : natural :=  666;      

	-- visable screen size in pixelsd
	constant X_VISIBLE : natural := 800; 
	constant Y_VISIBLE : natural := 600;
 
	constant FRAME_RATE : natural := 72;  -- frame rate in Hz
	constant VIDEO_LEN  : natural := 10;  -- video length in sec
	type matrix is array(natural range<>, natural range<>) of integer;
	constant jump : matrix(0 to 55, 0 to 48) :=(
		0=>(                           0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,12,12,12,12,12,9,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
		1=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,9,9,9,3,1,3,3,9,12,9,3,2,0,0,0,0,0,0,0,0,0,0,0,0),
		2=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,9,9,9,11,14,14,14,14,9,9,9,12,0,0,0,0,0,0,0,0,0,0,0,0),
		3=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,9,9,4,4,5,11,11,14,14,14,9,4,4,9,9,0,0,0,0,0,0,0,0,0,0,0),
		4=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,12,9,4,5,6,6,5,7,11,14,14,14,11,5,1,9,0,0,0,0,0,0,0,0,0,0,0),
		5=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,12,9,4,5,6,6,10,10,7,7,11,14,14,14,11,4,9,9,9,0,0,0,0,0,0,0,0,0),
		6=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,12,1,5,6,6,6,6,10,6,7,11,11,14,14,14,7,5,2,9,0,0,0,0,0,0,0,0,0),
		7=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,12,1,4,6,10,7,4,5,6,6,6,7,14,14,14,11,7,2,9,0,0,0,0,0,0,0,0,0),
		8=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,12,12,9,4,5,5,7,7,7,7,7,6,5,9,12,12,12,12,9,2,9,12,3,0,0,0,0,0,0,0),
		9=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,12,1,4,5,5,5,1,11,11,11,7,5,9,8,8,13,13,13,8,2,2,9,3,0,0,0,0,0,0,0),
	   10=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,12,1,1,1,1,5,11,11,11,11,11,11,5,9,8,12,15,13,13,2,1,9,3,0,0,0,0,0,0,0),
	   11=>(0,0,0,0,0,0,0,0,0,3,12,9,9,9,12,9,0,0,0,12,2,2,2,3,9,11,11,11,11,11,11,7,5,9,12,15,13,8,5,1,9,3,0,0,0,0,0,0,0),
	   12=>(0,0,0,0,0,0,0,0,0,9,9,2,2,2,3,12,0,0,0,12,2,2,3,12,12,1,11,11,1,1,1,11,11,5,8,13,4,7,11,5,9,3,0,0,0,0,0,0,0),
	   13=>(0,0,0,0,0,0,0,0,12,9,9,4,4,4,4,9,9,9,12,9,2,8,8,9,3,1,9,9,8,12,12,9,7,11,9,9,7,7,7,3,9,3,0,0,0,0,0,0,0),
	   14=>(0,0,0,0,0,0,3,9,12,1,5,5,5,5,5,1,1,3,1,1,2,8,13,3,2,2,8,8,8,12,15,9,5,11,7,7,11,7,2,3,9,3,0,0,0,0,0,0,0),
	   15=>(0,0,0,0,0,0,9,3,4,5,5,6,6,7,5,7,7,11,7,5,1,2,3,2,2,2,8,8,13,15,15,9,1,1,7,11,4,1,1,9,9,2,0,0,0,0,0,0,0),
	   16=>(0,0,0,0,0,12,9,4,4,5,6,6,6,6,5,11,11,14,11,11,1,4,5,1,4,4,9,8,13,15,15,9,3,9,12,11,1,9,9,9,0,0,0,0,0,0,0,0,0),
	   17=>(0,0,0,3,9,9,1,5,5,7,6,6,10,7,7,14,14,14,14,14,1,7,10,4,5,6,9,8,13,13,13,9,8,13,8,8,2,9,2,0,0,0,0,0,0,0,0,0,0),
	   18=>(0,0,0,9,12,12,9,5,6,6,6,10,10,6,7,14,14,14,14,11,1,7,10,4,4,5,9,8,13,13,13,13,13,13,13,13,3,9,2,0,0,0,0,0,0,0,0,0,0),
	   19=>(0,3,12,12,3,12,12,5,6,6,10,10,10,7,5,14,14,14,11,11,4,7,10,4,4,5,9,8,13,13,13,13,13,13,13,13,3,9,0,0,0,0,12,12,12,12,0,0,0),
	   20=>(0,9,9,9,12,15,15,15,14,7,6,6,5,4,1,3,3,3,1,4,10,6,6,4,4,5,5,9,15,13,8,3,8,13,13,8,2,9,0,0,0,2,12,3,3,12,3,0,0),
	   21=>(0,12,9,9,12,15,15,15,15,14,7,7,11,12,12,12,9,2,4,5,7,7,5,4,4,5,7,5,12,13,13,12,8,13,8,9,12,12,0,0,12,12,9,9,9,9,12,9,0),
	   22=>(0,12,9,9,12,15,15,15,15,15,9,9,9,0,2,2,9,3,4,5,5,4,1,5,5,7,6,6,9,12,12,12,12,8,3,9,12,0,0,9,12,3,9,12,12,12,3,12,9),
	   23=>(0,12,9,9,12,15,15,15,15,15,9,9,9,0,0,0,9,12,9,1,1,4,5,5,7,6,6,10,6,7,9,9,9,3,12,12,3,0,3,12,9,12,9,3,12,12,12,9,9),
	   24=>(0,9,12,9,12,15,15,15,15,15,12,12,9,0,0,0,0,3,9,1,9,4,4,5,6,6,10,10,6,6,7,5,4,4,12,9,9,9,9,9,4,12,9,3,12,12,12,9,9),
	   25=>(0,0,3,9,2,12,12,12,9,3,12,3,0,0,0,0,0,3,9,4,11,7,1,5,6,6,10,10,10,10,10,5,4,7,4,3,12,9,1,4,5,1,2,3,12,12,12,9,9),
	   26=>(0,0,0,9,9,9,9,9,9,9,9,0,0,0,0,0,9,9,9,7,14,11,7,4,5,6,6,6,10,10,6,4,4,7,7,5,9,9,4,5,5,9,12,9,9,9,12,9,9),
	   27=>(0,0,0,0,0,9,3,3,12,0,0,0,0,0,0,0,9,1,5,7,14,14,11,3,1,5,7,6,10,6,6,4,4,7,7,7,4,4,5,5,5,12,12,12,3,9,12,9,9),
	   28=>(0,0,0,0,0,3,3,3,3,0,0,0,0,0,0,0,9,2,1,1,3,3,3,2,2,1,4,4,5,5,4,7,7,7,7,7,5,5,5,5,5,3,9,12,12,9,3,12,3),
	   29=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,1,1,4,5,5,7,7,12,12,7,5,4,1,1,12,14,5,7,7,5,5,5,5,5,4,9,9,12,9,2,12,0),
	   30=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,1,4,5,7,11,11,14,14,14,14,11,4,1,3,15,15,3,5,7,4,4,5,5,5,5,4,2,2,2,2,12,0),
	   31=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,2,4,7,14,14,14,14,14,14,12,7,7,6,7,9,12,15,9,4,4,5,5,5,5,1,1,3,12,12,12,9,0),
	   32=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,9,9,2,4,7,14,14,14,14,14,14,9,4,10,10,6,5,9,12,12,9,4,5,5,4,4,9,9,9,9,0,0,0,0),
	   33=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,3,1,2,4,7,11,14,14,11,11,7,4,4,11,10,10,10,7,3,12,15,3,1,1,2,9,9,9,9,3,0,0,0,0),
	   34=>(0,0,0,0,0,0,0,0,12,9,9,9,9,9,9,5,7,7,5,4,7,7,7,7,7,5,4,5,10,10,10,10,10,7,12,12,12,12,12,12,12,3,0,0,0,0,0,0,0),
	   35=>(0,2,9,9,9,9,9,9,12,2,2,1,2,2,1,7,11,11,5,1,1,1,2,2,2,1,4,5,10,10,10,10,10,10,5,9,12,9,9,9,9,9,9,9,9,9,0,0,0),
	   36=>(0,9,9,9,9,9,9,9,4,5,5,5,5,4,1,7,11,11,11,11,7,4,3,12,9,1,4,5,10,10,10,10,10,10,6,6,9,9,9,9,9,9,9,9,9,12,9,0,0),
	   37=>(12,12,9,1,1,1,1,4,5,5,5,5,5,4,4,5,7,11,11,11,5,9,12,12,9,1,4,7,10,10,10,10,10,10,6,6,4,4,5,5,5,5,5,5,5,9,12,9,0),
	   38=>(12,1,5,4,1,4,5,5,5,5,5,5,5,5,5,1,7,11,7,7,1,9,0,0,9,1,4,6,6,6,10,10,10,10,6,6,4,7,10,10,10,10,10,10,10,7,1,12,0),
	   39=>(12,1,5,4,1,4,5,5,5,5,5,5,7,7,7,4,5,7,4,9,9,12,0,0,9,1,4,5,7,6,10,10,10,10,7,5,7,6,10,10,10,10,10,6,5,4,2,12,0),
	   40=>(12,1,5,4,1,4,5,5,5,5,5,5,7,7,7,5,5,1,2,9,3,0,0,0,9,9,4,5,5,6,10,10,10,10,5,4,6,6,10,10,10,10,6,6,4,3,3,12,0),
	   41=>(12,1,5,4,1,4,5,5,5,7,7,7,7,7,7,7,7,5,1,9,3,0,0,0,9,9,9,4,5,6,6,10,10,10,5,4,10,10,10,10,10,6,5,1,1,12,12,3,0),
	   42=>(12,1,5,5,4,4,5,5,5,7,7,7,7,7,7,7,5,4,9,12,3,0,0,0,0,0,9,1,5,7,6,6,6,6,5,4,10,10,10,10,6,7,4,3,12,12,3,0,0),
	   43=>(12,1,5,5,5,4,4,5,5,7,7,7,7,7,7,5,4,1,9,0,0,0,0,0,0,0,9,1,4,5,7,6,6,6,5,4,10,10,10,6,6,1,1,3,9,0,0,0,0),
	   44=>(12,1,5,5,7,5,4,4,5,5,7,7,5,4,4,1,9,12,9,0,0,0,0,0,0,0,12,12,3,4,5,6,7,5,7,6,10,10,6,5,4,1,9,12,9,0,0,0,0),
	   45=>(12,1,5,5,7,7,5,4,4,4,5,5,4,9,9,9,9,0,0,0,0,0,0,0,0,0,0,9,9,9,4,4,4,4,7,6,10,6,6,4,3,9,9,0,0,0,0,0,0),
	   46=>(12,1,5,5,7,7,7,5,4,1,1,1,1,12,3,9,2,0,0,0,0,0,0,0,0,0,0,0,2,12,1,1,4,5,5,7,6,7,4,1,9,9,3,0,0,0,0,0,0),
	   47=>(9,9,3,4,7,7,7,7,5,4,1,9,9,9,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,9,9,1,5,5,5,5,4,1,9,9,3,0,0,0,0,0,0,0),
	   48=>(0,12,9,4,7,7,7,7,7,5,1,9,9,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,9,1,5,5,5,1,1,3,9,0,0,0,0,0,0,0,0,0),
	   49=>(0,12,9,1,5,7,7,7,7,5,1,9,9,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,9,4,5,5,5,1,9,9,3,0,0,0,0,0,0,0,0,0),
	   50=>(0,9,12,9,4,7,7,7,5,4,9,12,9,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,12,9,4,4,4,12,12,0,0,0,0,0,0,0,0,0,0,0),
	   51=>(0,0,2,9,1,5,7,7,5,3,12,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,12,3,1,3,12,2,0,0,0,0,0,0,0,0,0,0,0),
	   52=>(0,0,0,9,1,5,7,5,4,3,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,12,12,12,9,0,0,0,0,0,0,0,0,0,0,0,0),
	   53=>(0,0,0,9,9,5,7,5,4,9,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	   54=>(0,0,0,9,12,9,1,1,12,12,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	   55=>(0,0,0,0,0,12,12,12,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0)
	   
	);
	constant still : matrix(0 to 55, 0 to 48) :=(
		0=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,12,12,9,9,9,9,9,9,12,0,0,0,0,0,0,0,0,0,0,0,0),
		1=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,9,9,9,12,9,4,9,9,9,9,9,12,9,9,9,9,9,0,0,0,0,0,0,0),
		2=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,9,2,2,2,3,14,11,14,14,14,14,14,9,1,2,2,3,9,0,0,0,0,0,0,0),
		3=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,9,9,9,4,4,4,5,7,11,11,11,11,14,14,14,12,11,11,6,9,9,9,0,0,0,0,0),
		4=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,9,12,1,1,4,5,5,5,6,7,7,5,4,4,11,11,14,14,14,14,11,4,1,9,12,9,3,0,0),
		5=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,12,9,9,4,5,5,5,6,7,7,10,10,7,7,6,4,4,5,11,11,14,14,6,5,4,9,9,12,0,0),
		6=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,2,4,5,5,6,6,7,7,7,7,10,7,7,6,5,5,5,5,11,14,14,11,11,5,1,9,12,0,0),
		7=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,1,4,5,6,7,7,7,7,7,6,6,5,5,6,7,7,5,1,9,14,14,14,14,12,2,9,12,0,0),
		8=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,12,12,12,9,4,5,5,6,7,7,7,6,5,11,11,11,11,11,6,6,4,8,9,12,12,13,12,9,8,8,12,12,12),
		9=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,3,1,4,5,5,5,5,6,6,5,4,4,11,11,11,11,11,5,5,9,8,8,13,13,13,13,13,8,8,2,2,12),
	   10=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,3,1,4,5,4,4,4,4,4,5,11,11,11,11,11,11,11,11,11,5,5,9,8,8,15,15,12,8,8,2,2,12),
	   11=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,3,1,4,4,4,1,1,9,9,9,11,11,11,11,11,11,11,11,11,6,6,5,9,9,12,15,12,9,3,1,2,12),
	   12=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,3,2,1,1,2,2,2,12,12,9,2,1,14,11,5,1,2,1,1,11,11,11,5,5,8,13,8,4,4,1,2,12),
	   13=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,3,2,2,2,3,8,8,8,9,3,2,2,9,9,9,8,12,15,15,9,5,5,11,11,5,9,5,11,11,1,2,12),
	   14=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,9,9,9,3,2,8,13,13,8,2,2,2,2,8,8,8,13,12,15,15,9,1,4,14,11,5,5,11,11,14,9,9,12),
	   15=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,3,9,9,9,2,8,13,13,8,2,2,2,2,8,8,13,13,15,15,15,9,2,1,1,4,11,10,5,1,9,12,9,3),
	   16=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,12,12,12,12,14,6,5,5,9,9,3,2,2,3,8,8,8,13,13,13,15,15,9,2,9,12,12,5,6,9,9,12,9,0,0),
	   17=>(0,0,0,0,0,0,0,0,0,0,0,0,9,12,12,1,1,4,5,6,7,7,10,11,5,1,3,8,8,8,8,13,13,13,13,13,8,2,9,13,13,3,3,9,0,0,0,0,0),
	   18=>(0,0,0,0,0,0,0,0,0,0,0,12,12,9,9,2,1,1,4,4,4,5,7,7,7,11,5,3,3,8,8,13,13,13,13,13,13,13,13,13,13,12,9,12,0,0,0,0,0),
	   19=>(0,0,0,0,0,0,0,0,0,0,0,12,12,2,1,4,4,5,5,4,4,5,6,6,10,10,6,1,2,8,8,13,13,13,13,13,13,13,13,13,13,12,12,12,0,0,0,0,0),
	   20=>(0,0,0,0,0,0,0,0,0,0,0,12,12,1,4,5,6,11,11,11,5,5,4,4,11,10,6,1,2,8,8,13,13,13,3,2,13,13,13,13,13,3,3,9,0,0,0,0,0),
	   21=>(0,0,0,0,0,0,0,0,0,12,12,12,9,5,6,11,11,14,14,14,11,11,1,4,6,7,5,1,2,3,3,8,13,13,13,13,13,13,13,8,9,12,12,12,0,0,0,0,0),
	   22=>(0,0,0,0,0,0,0,3,3,12,3,1,5,5,11,11,11,14,14,14,11,11,1,4,6,7,5,4,1,1,2,8,8,8,13,13,13,13,8,3,3,9,0,0,0,0,0,0,0),
	   23=>(0,0,0,0,0,0,2,12,9,9,4,5,5,6,5,5,6,14,14,14,6,5,1,1,1,4,5,11,11,4,1,2,2,2,3,3,3,3,9,12,9,3,0,0,0,0,0,0,0),
	   24=>(0,0,0,0,0,0,0,9,2,1,5,5,6,6,6,6,6,11,14,11,5,4,1,1,2,1,5,11,11,4,1,2,2,3,9,9,9,9,9,0,0,0,0,0,0,0,0,0,0),
	   25=>(0,0,0,0,0,0,0,3,2,1,5,5,7,10,10,10,10,6,5,4,1,1,1,1,1,1,5,11,11,4,1,1,1,9,12,2,2,2,2,0,0,0,0,0,0,0,0,0,0),
	   26=>(0,0,0,0,0,0,0,3,2,1,5,6,7,7,7,10,10,6,6,5,4,4,12,12,12,12,12,5,5,4,4,5,6,5,12,12,12,12,12,0,0,0,0,0,0,0,0,0,0),
	   27=>(0,0,0,0,0,0,0,9,9,9,4,5,6,7,7,10,10,7,7,6,5,9,12,12,15,15,12,9,3,4,5,6,7,11,3,3,3,3,9,12,12,9,0,0,0,0,0,0,0),
	   28=>(0,0,0,0,0,0,0,9,12,12,3,1,5,6,6,7,7,7,5,11,12,12,15,15,15,15,15,15,15,9,1,1,4,3,12,12,12,12,12,3,9,9,0,0,0,0,0,0,0),
	   29=>(0,0,0,0,0,0,0,0,0,12,3,1,4,6,6,6,6,6,5,12,12,15,15,15,15,15,15,15,15,9,2,3,9,9,9,9,9,9,9,9,9,9,9,12,0,0,0,0,0),
	   30=>(0,0,0,0,0,0,0,0,0,12,3,2,4,6,5,5,5,5,5,12,12,15,15,15,15,15,15,15,15,9,2,9,12,12,3,2,2,2,9,12,12,3,2,9,0,0,0,0,0),
	   31=>(0,0,0,0,0,0,0,0,0,12,3,1,6,11,11,4,4,5,5,12,12,15,15,15,15,15,15,15,15,9,2,9,12,12,3,2,9,12,12,12,12,3,2,9,0,0,0,0,0),
	   32=>(0,0,0,0,0,0,0,0,0,12,3,1,11,11,11,9,9,4,4,9,12,12,15,15,15,15,15,15,15,9,9,9,12,9,9,9,12,12,12,12,12,9,9,12,0,0,0,0,0),
	   33=>(0,0,0,0,0,0,0,0,0,12,3,1,6,11,14,14,14,3,1,1,2,9,12,12,12,12,12,3,3,12,12,12,2,3,12,12,12,12,12,2,3,12,12,9,0,0,0,0,0),
	   34=>(0,0,0,0,0,0,2,12,12,12,2,1,6,11,14,14,14,14,11,5,4,4,9,9,9,9,9,2,3,12,2,12,12,12,9,9,9,9,9,12,12,9,0,0,0,0,0,0,0),
	   35=>(0,0,0,0,0,12,12,9,1,1,1,1,4,5,11,14,14,14,14,14,6,5,1,1,1,1,1,2,3,12,0,0,0,12,9,3,3,3,9,0,0,0,0,0,0,0,0,0,0),
	   36=>(0,0,0,0,12,9,9,4,5,5,4,4,4,4,11,14,14,14,14,14,11,11,1,1,11,14,9,1,3,12,0,0,0,9,12,9,9,9,12,0,0,0,0,0,0,0,0,0,0),
	   37=>(0,0,12,12,12,4,4,4,5,5,5,5,4,1,4,11,11,14,14,14,14,9,1,1,14,11,11,4,4,12,12,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	   38=>(0,0,12,2,1,4,5,5,5,5,5,5,4,1,4,5,5,4,1,1,1,1,2,1,11,11,11,5,5,1,1,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	   39=>(0,0,12,2,1,5,5,5,5,5,4,4,4,4,5,5,5,6,6,6,6,5,1,1,5,11,6,5,5,4,1,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	   40=>(12,12,12,3,4,5,5,5,5,4,1,4,5,6,6,5,6,7,7,10,10,11,4,1,4,5,5,5,5,4,1,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	   41=>(12,9,4,5,5,5,5,4,1,1,5,5,6,7,7,10,10,10,10,10,10,11,1,1,4,5,5,5,5,4,2,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	   42=>(9,2,4,5,5,5,4,4,4,5,6,6,7,7,10,10,10,10,10,10,10,11,4,1,4,5,5,5,4,1,2,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	   43=>(9,1,4,5,5,1,1,4,5,6,7,7,10,10,10,10,10,10,10,10,10,11,4,1,4,5,5,5,4,1,2,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	   44=>(9,1,4,5,5,1,1,4,5,6,7,7,10,10,10,10,10,10,10,10,10,11,4,1,1,4,4,4,4,12,12,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	   45=>(12,9,4,5,5,1,1,4,5,6,7,7,10,10,10,10,10,10,10,10,10,6,4,2,3,9,9,9,9,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	   46=>(3,2,12,3,1,2,1,4,5,6,7,7,10,10,10,10,10,10,10,10,7,6,4,2,12,3,3,3,3,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	   47=>(0,0,12,9,9,3,2,4,5,6,7,7,10,10,10,10,10,10,10,6,6,5,4,2,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	   48=>(0,0,0,0,12,3,2,4,5,6,7,7,10,10,10,10,10,7,6,5,4,1,1,1,12,9,9,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	   49=>(0,0,0,0,12,9,1,4,5,5,6,6,7,7,7,7,7,5,5,5,11,7,6,6,9,9,12,3,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	   50=>(0,0,12,12,12,4,4,4,4,4,5,5,6,6,6,6,6,5,4,11,10,10,7,7,6,4,9,12,12,9,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	   51=>(0,0,12,3,1,5,5,4,1,1,1,1,1,4,4,1,4,11,10,10,10,10,10,10,7,7,5,4,3,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	   52=>(0,0,12,2,1,5,5,5,4,4,4,4,5,6,5,6,6,10,10,10,10,10,10,10,10,10,7,6,5,9,9,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	   53=>(0,0,12,2,1,4,5,5,5,5,5,5,6,7,7,11,10,10,10,10,10,11,11,10,10,10,10,7,6,4,1,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	   54=>(0,0,12,2,1,1,1,1,1,1,1,1,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,1,1,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
	   55=>(0,0,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0)
	);
constant run : matrix(0 to 55, 0 to 48) :=(
	0=>(                                     0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,12,8,8,8,8,12,0,0,0,0,0,0,0,0,0,0,0,0,0),
	1=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,8,8,8,8,3,2,2,2,12,8,8,8,2,0,0,0,0,0,0,0,0,0),
	2=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,12,8,1,1,9,13,13,13,13,12,1,1,8,8,0,0,0,0,0,0,0,0,0),
	3=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,12,12,8,3,3,9,10,13,13,13,13,9,9,8,12,12,0,0,0,0,0,0,0,0),
	4=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,2,8,8,1,4,4,4,6,5,3,8,13,13,13,13,13,1,12,8,2,0,0,0,0,0,0),
	5=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8,8,8,3,4,4,6,6,10,9,9,3,9,9,13,13,4,8,8,12,0,0,0,0,0,0),
	6=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8,1,3,4,4,6,5,6,10,10,9,3,4,9,13,13,9,3,2,12,0,0,0,0,0,0),
	7=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8,1,3,4,5,5,10,9,4,4,6,6,4,2,13,13,13,8,1,12,0,0,0,0,0,0),
	8=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8,12,8,3,4,4,5,5,9,9,9,9,9,6,4,2,12,12,12,8,8,12,12,2,0,0,0,0),
	9=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8,8,1,4,4,4,6,6,2,9,13,10,10,4,8,7,11,11,11,11,7,1,8,8,0,0,0,0),
   10=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8,8,1,4,3,3,3,4,13,10,10,13,10,10,9,8,7,11,14,11,7,2,8,8,0,0,0,0),
   11=>(0,0,0,0,0,0,0,0,0,0,0,0,0,2,8,8,8,8,8,0,0,8,8,1,3,2,1,1,8,13,13,13,13,13,13,9,4,8,12,15,12,8,2,8,8,0,0,0,0),
   12=>(0,0,0,0,0,0,0,0,0,0,0,0,0,8,2,2,2,2,12,2,0,8,8,1,1,1,1,12,12,1,9,13,3,1,1,9,10,4,8,11,8,3,1,8,8,0,0,0,0),
   13=>(0,0,0,0,0,0,0,0,0,0,0,8,12,12,2,3,3,3,8,12,12,12,2,1,1,7,7,8,8,1,8,12,8,8,12,12,9,9,4,7,8,9,2,8,8,0,0,0,0),
   14=>(0,0,0,0,0,0,0,0,0,0,2,8,2,3,3,4,4,4,3,1,1,1,1,1,0,7,11,2,0,0,2,7,7,12,15,12,1,13,10,4,9,13,2,8,8,0,0,0,0),
   15=>(0,0,0,0,0,0,0,0,0,0,12,12,3,4,4,6,6,4,4,4,9,9,4,3,1,2,7,1,0,0,7,7,11,14,15,12,1,8,9,9,9,8,12,8,2,0,0,0,0),
   16=>(0,0,0,0,0,0,0,0,8,12,8,2,4,4,6,6,5,6,4,9,13,13,9,9,1,1,2,1,1,1,7,7,14,14,15,12,0,2,3,9,4,2,12,0,0,0,0,0,0),
   17=>(0,0,0,0,0,0,0,0,12,2,3,4,4,6,5,6,10,9,9,13,13,13,13,13,1,4,9,2,3,9,8,7,14,14,14,12,1,12,12,2,12,8,8,0,0,0,0,0,0),
   18=>(0,0,0,0,0,0,8,12,12,8,3,4,6,6,6,10,10,9,9,13,13,13,13,13,1,9,10,2,1,4,8,7,14,14,14,11,7,14,14,12,12,0,0,0,0,0,0,0,0),
   19=>(0,0,0,0,0,1,12,8,8,12,8,4,5,5,10,10,10,4,9,13,13,13,13,13,1,9,10,2,0,1,2,7,14,14,14,14,14,11,12,12,2,0,0,0,0,0,0,0,0),
   20=>(0,0,0,0,0,12,12,12,12,15,15,13,9,6,10,10,9,3,3,8,8,8,8,9,6,9,10,3,0,0,7,7,14,14,7,11,14,14,14,12,12,0,0,0,0,0,0,0,0),
   21=>(0,0,0,0,0,12,1,12,12,15,15,15,8,9,10,9,3,2,2,0,0,1,1,3,5,6,10,3,1,1,7,7,14,11,2,11,14,14,14,2,12,1,2,2,2,2,0,0,0),
   22=>(0,0,0,0,0,12,1,12,12,15,15,15,15,12,1,12,15,15,12,1,1,1,3,9,10,9,3,3,4,10,4,2,7,11,14,14,11,7,8,12,8,8,8,8,8,12,0,0,0),
   23=>(0,0,0,0,0,12,1,12,12,15,15,15,15,12,1,12,15,15,15,1,3,8,3,4,9,4,3,4,9,10,9,3,8,7,11,11,7,8,8,8,8,8,8,8,8,12,8,8,0),
   24=>(0,0,0,0,0,12,2,12,12,15,15,15,15,12,1,12,15,15,15,1,9,13,2,1,1,3,4,10,10,10,6,6,3,1,0,1,1,12,0,0,12,1,12,12,12,8,1,8,0),
   25=>(0,0,0,0,0,8,12,8,12,15,15,15,12,12,12,15,15,12,12,3,9,13,13,8,1,4,6,10,10,10,5,5,3,1,4,3,1,12,12,12,8,8,8,8,12,12,8,12,12),
   26=>(0,0,0,0,0,0,12,8,2,12,12,12,2,12,15,15,15,8,3,3,9,10,13,13,2,4,5,6,10,10,6,6,3,3,9,4,2,12,12,1,8,12,2,2,12,12,12,2,8),
   27=>(0,0,0,0,0,0,12,8,1,2,2,2,15,15,15,12,8,3,4,4,4,9,13,13,13,9,4,6,5,6,6,3,9,10,10,9,4,8,8,1,8,12,2,2,12,12,12,2,8),
   28=>(0,0,0,0,0,8,12,8,1,1,2,2,12,15,15,12,1,4,4,4,4,4,13,13,13,9,3,6,6,6,4,1,9,10,10,10,9,3,1,2,8,12,8,8,12,12,12,2,8),
   29=>(0,0,0,0,2,12,2,3,4,4,4,3,1,12,15,12,1,4,4,4,4,4,2,9,13,13,9,3,1,1,1,1,4,9,10,13,13,3,3,4,6,6,12,12,1,8,12,2,8),
   30=>(0,0,0,8,8,8,3,4,4,3,3,3,3,8,12,8,1,4,4,4,9,9,13,12,9,8,3,12,12,12,12,12,8,4,9,9,9,3,4,6,5,5,9,9,8,8,8,2,8),
   31=>(0,0,0,8,1,3,4,4,3,1,1,3,3,3,2,1,1,3,4,4,9,13,13,13,1,1,1,8,0,0,0,2,8,3,9,3,1,4,6,5,5,5,5,6,12,8,1,1,8),
   32=>(0,0,0,8,1,3,4,3,3,3,4,3,4,4,3,3,1,1,3,9,13,13,13,13,13,8,1,8,0,0,0,2,12,12,2,1,1,6,5,5,5,5,6,4,2,1,1,12,12),
   33=>(0,1,12,8,2,4,4,1,2,4,4,4,4,4,4,3,1,1,2,9,13,13,13,13,13,9,2,12,12,0,0,0,0,8,8,2,1,6,5,5,5,5,4,3,8,8,8,8,0),
   34=>(0,2,8,2,4,6,6,3,2,4,4,4,4,4,4,4,3,1,3,9,9,13,13,13,13,13,9,3,8,8,0,0,0,2,8,8,1,4,4,4,4,4,3,8,8,8,8,2,0),
   35=>(0,2,8,3,6,5,5,3,2,4,4,6,6,6,4,3,3,3,3,4,9,9,13,13,13,13,4,4,9,12,12,0,0,0,0,12,12,8,3,3,3,3,12,12,8,0,0,0,0),
   36=>(8,12,8,4,5,5,5,4,3,4,6,5,5,6,4,3,2,9,4,2,4,9,10,13,13,9,1,6,6,3,12,8,2,0,0,0,8,8,1,1,1,2,12,0,0,0,0,0,0),
   37=>(12,8,3,6,5,5,5,6,4,3,4,6,5,5,5,4,1,9,9,13,8,3,9,9,13,9,1,9,6,6,4,8,12,0,0,0,1,12,12,12,12,12,8,0,0,0,0,0,0),
   38=>(12,1,4,6,5,5,5,5,6,3,3,4,6,5,5,6,3,4,9,13,9,3,4,9,13,9,4,10,10,5,4,1,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
   39=>(12,1,6,5,5,5,5,5,6,4,3,3,4,6,5,5,6,3,4,13,9,9,3,1,1,4,5,10,10,10,9,2,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
   40=>(12,2,6,5,5,5,5,6,4,3,8,12,2,3,4,5,6,3,3,10,9,4,1,1,3,9,6,10,10,10,9,4,12,12,2,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
   41=>(12,1,6,5,5,5,5,4,3,1,12,2,8,1,1,4,6,3,2,9,3,1,0,1,4,9,10,10,10,10,6,6,3,8,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
   42=>(12,1,6,5,6,4,3,3,8,12,12,2,12,12,12,12,3,1,1,2,12,12,8,2,4,9,10,10,10,10,10,10,3,8,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
   43=>(12,8,6,6,4,3,8,8,12,8,0,0,0,0,2,12,8,8,8,8,12,8,8,1,4,9,10,10,10,10,10,10,3,8,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
   44=>(2,8,8,1,1,8,8,8,8,0,0,0,0,0,0,2,8,8,8,8,2,8,8,1,4,9,10,10,10,10,10,10,3,8,12,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
   45=>(0,2,8,8,8,8,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8,8,1,4,6,10,10,10,10,10,9,1,8,12,8,0,0,0,0,0,0,0,0,0,0,0,0,0),
   46=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8,8,2,4,6,5,10,10,10,9,1,1,1,1,12,8,8,2,0,0,0,0,0,0,0,0,0,0),
   47=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8,8,2,4,4,6,6,6,4,4,6,9,9,6,8,12,12,12,2,0,0,0,0,0,0,0,0,0),
   48=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8,8,1,4,4,4,6,6,3,4,5,10,10,6,6,3,2,8,12,8,0,0,0,0,0,0,0,0),
   49=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8,8,1,4,4,4,3,3,6,6,10,10,10,10,10,10,6,9,8,12,0,0,0,0,0,0,0,0),
   50=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8,12,8,3,3,3,3,4,6,10,10,10,10,10,10,10,6,6,4,8,8,8,0,0,0,0,0,0),
   51=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8,12,1,1,1,4,4,10,10,10,10,10,10,10,10,10,10,6,4,2,12,0,0,0,0,0,0),
   52=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8,1,1,3,4,4,6,10,10,10,10,10,10,6,6,9,4,3,2,12,0,0,0,0,0,0),
   53=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8,2,3,4,4,4,6,6,10,10,10,10,6,6,4,3,2,2,2,12,0,0,0,0,0,0),
   54=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8,12,12,1,1,1,3,3,3,3,3,3,3,3,2,8,12,12,12,1,0,0,0,0,0,0),
   55=>(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8,12,12,12,12,12,12,12,12,12,12,12,12,12,2,0,0,0,0,0,0,0,0,0)   
	);
-- spiral demo constants -------------------------------
type RAM is array(natural range<>) of integer;
	signal LUT : RAM(0 to 15) := (16#000000#, 16#0000AA#, 16#00AA00#, 16#00AAAA#, 16#AA0000#, 16#AA00AA#, 16#AA5500#, 16#AAAAAA#, 16#555555#, 16#5555ff#, 16#55ff55#, 16#55ffff#, 16#ff5555#,16#ff55ff#,16#ffff55#,16#ffffff#);
	--type pixel is integer;

	constant STEP_WIDTH : natural := 32;
	constant X_START : natural :=  325;  
	signal Y_START : natural := 296;   

-- spiral demo signals ---------------------------------
-- registers
	-- states
	-- states
	type state_t is (drawPixel,updateBitMap);
	type image_t is (run_s, jump_s, still_s);
	signal state, stateNext : state_t := (drawPixel);
	-- temp. video stream for assembling components  
	signal videoStreamOutTemp, videoStreamOutTempNext : VideoStream_t := VIDEO_STREAM_IDLE;
	-- current upper right corner of square
	constant imageWidth : natural := 48;
	constant imageHeight : natural := 55;
	signal currentPixelY : natural range 0 to 55;
	signal frameCounter : natural range 0 to 10;
	signal pixelHoldX : natural range 0 to 6;
	signal pixelHoldY : natural range 0 to 6;
	signal currentMap : matrix(0 to 55, 0 to 48);
	signal currentImage : image_t;
	signal nextImage: image_t;
	signal xPos : natural range 0 to X_FULL-1 := 0; 
	signal yPos : natural range 0 to Y_FULL-1 := 0; 
	signal currentColour : integer range 0 to 16777215;
	signal jumpCounter : natural range 0 to 5;
	signal doWhile : std_logic := '1';

	signal jumpConditionMet : std_logic := '0';
begin

-- forward video stream register to output 
videoStreamOut <= videoStreamOutTemp; 


-- sequential process with registers
reset : process (clk)
variable previousY : natural range 1 to Y_FULL-1;
variable currentPixelX : natural range 0 to 48;
begin

	if rising_edge(clk) then    
		if sresetn = '0' then
			state 			<= drawPixel 	after 2 ns; 
			jumpConditionMet 	<= '0';
			currentImage <= still_s;
			frameCounter <= 0;
			currentPixelX := 0;
			pixelHoldY <= 0;
			currentMap <= still;
			videoStreamOutTemp <= VIDEO_STREAM_IDLE after 2 ns;
			previousY := Y_START;
			currentColour <= 0;
			jumpCounter <= 0;
			doWhile <= '1';
		else
			state <= stateNext 			after 2 ns;
			currentImage <= nextImage; 
			videoStreamOutTemp <= videoStreamOutTempNext after 2 ns;
			yPos <= to_integer(videoStreamIn.verticalPos);  			-- rename current x,y position for easier handling 
			xPos <= to_integer(videoStreamIn.horizontalPos);
			videoStreamOutTempNext <= videoStreamIn after 2 ns; 		-- copy input video stream to temp register                     
			if AUDIO_IN(W - 2) = '1' then -- audio in not yet implemented
				jumpConditionMet <= '1';  
			end if;
				case state is
					when drawPixel 	=> 
					if(not((yPos >= Y_START and yPos < (Y_START + (imageHeight * 4))) and (xPos >= X_START and (xPos < (X_START + (imageWidth * 4)))))) then
							if(yPos = (Y_FULL - 10)) then
								currentPixelY <= 0;
								previousY := Y_START;
							end if;
							if(xPos = (X_FULL - 1)) then
								currentPixelX := 0;
							end if;
							if(yPos > X_START + (4 * imageWidth)) then
								videoStreamOutTempNext.pixelRGBData <= to_unsigned(6697728,NUM_BITS_PIXEL_RGB);
							else
								videoStreamOutTempNext.pixelRGBData <= to_unsigned(0,NUM_BITS_PIXEL_RGB);
							end if;
					else
							if doWhile = '1' then 
								currentColour <= LUT(currentMap(currentPixelY, currentPixelX));
								doWhile <= '0';
							end if;
							if pixelHoldX = 3 then
							pixelHoldX <= 0;
							currentPixelX := currentPixelX + 1;
							doWhile <= '1';
						else
							pixelHoldX <= pixelHoldX + 1;
						end if;
						if((yPos - previousY) = 4) then
							previousY := yPos;
							doWhile <= '1';
							currentPixelY <= currentPixelY + 1;
						end if;
						videoStreamOutTempNext.pixelRGBData <= to_unsigned(currentColour, NUM_BITS_PIXEL_RGB);
					end if;
					if (yPos = (Y_FULL - 1) and xPos = (X_FULL - 1)) then
						stateNext <= updateBitMap; 
					end if;
					when updateBitMap  =>
						stateNext <= drawPixel;
						if frameCounter = 1 then
							frameCounter <= 0;
							if jumpConditionMet = '1' then							
								if jumpCounter = 0 then
								jumpCounter <= jumpCounter + 1;
								currentMap <= jump;
								currentImage <= jump_s;
								Y_START <= 225;
								previousY := 225;
								elsif jumpCounter = 1 then
									Y_START <= 200;
									previousY := 200;
									jumpCounter <= jumpCounter + 1;
									
								elsif jumpCounter = 2 then
									Y_START <= 225;
									previousY := 225;
									jumpCounter <= jumpCounter + 1;
								elsif jumpCounter = 3 then
									Y_START <= 296;
									previousY := 296;
									jumpCounter <= 0;
									nextImage <= still_s;
									jumpConditionMet <= '0'; 
								end if;
							elsif currentImage = jump_s then 
								currentMap <= still;
								nextImage <= still_s;			
							elsif currentImage = run_s then
								currentMap <= still;
								nextImage <= still_s;
							elsif currentImage = still_s then
								currentMap <= run;
								nextImage <= run_s;
							end if;
						else
							frameCounter <= frameCounter + 1;
						end if;

				end case;
		end if;
	end if;
end process;


end architecture RTL;


